
module InvSubBytes(stateIn,stateOut);


input wire[127:0] stateIn;
output wire[127:0] stateOut;

    
wire [2047:0] c;



assign  c[7:0]=8'h52;
assign  c[15:8]=8'h09;
assign  c[23:16]=8'h6a;
assign  c[31:24]=8'hd5;
assign  c[39:32]=8'h30;
assign  c[47:40]=8'h36;
assign  c[55:48]=8'ha5;
assign  c[63:56]=8'h38;
assign  c[71:64]=8'hbf;
assign  c[79:72]=8'h40;
assign  c[87:80]=8'ha3;
assign  c[95:88]=8'h9e;
assign  c[103:96]=8'h81;
assign  c[111:104]=8'hf3;
assign  c[119:112]=8'hd7;
assign  c[127:120]=8'hfb;
assign  c[135:128]=8'h7c;
assign  c[143:136]=8'he3;
assign  c[151:144]=8'h39;
assign  c[159:152]=8'h82;
assign  c[167:160]=8'h9b;
assign  c[175:168]=8'h2f;
assign  c[183:176]=8'hff;
assign  c[191:184]=8'h87;
assign  c[199:192]=8'h34;
assign  c[207:200]=8'h8e;
assign  c[215:208]=8'h43;
assign  c[223:216]=8'h44;
assign  c[231:224]=8'hc4;
assign  c[239:232]=8'hde;
assign  c[247:240]=8'he9;
assign  c[255:248]=8'hcb;
assign  c[263:256]=8'h54;
assign  c[271:264]=8'h7b;
assign  c[279:272]=8'h94;
assign  c[287:280]=8'h32;
assign  c[295:288]=8'ha6;
assign  c[303:296]=8'hc2;
assign  c[311:304]=8'h23;
assign  c[319:312]=8'h3d;
assign  c[327:320]=8'hee;
assign  c[335:328]=8'h4c;
assign  c[343:336]=8'h95;
assign  c[351:344]=8'h0b;
assign  c[359:352]=8'h42;
assign  c[367:360]=8'hfa;
assign  c[375:368]=8'hc3;
assign  c[383:376]=8'h4e;
assign  c[391:384]=8'h08;
assign  c[399:392]=8'h2e;
assign  c[407:400]=8'ha1;
assign  c[415:408]=8'h66;
assign  c[423:416]=8'h28;
assign  c[431:424]=8'hd9;
assign  c[439:432]=8'h24;
assign  c[447:440]=8'hb2;
assign  c[455:448]=8'h76;
assign  c[463:456]=8'h5b;
assign  c[471:464]=8'ha2;
assign  c[479:472]=8'h49;
assign  c[487:480]=8'h6d;
assign  c[495:488]=8'h8b;
assign  c[503:496]=8'hd1;
assign  c[511:504]=8'h25;
assign  c[519:512]=8'h72;
assign  c[527:520]=8'hf8;
assign  c[535:528]=8'hf6;
assign  c[543:536]=8'h64;
assign  c[551:544]=8'h86;
assign  c[559:552]=8'h68;
assign  c[567:560]=8'h98;
assign  c[575:568]=8'h16;
assign  c[583:576]=8'hd4;
assign  c[591:584]=8'ha4;
assign  c[599:592]=8'h5c;
assign  c[607:600]=8'hcc;
assign  c[615:608]=8'h5d;
assign  c[623:616]=8'h65;
assign  c[631:624]=8'hb6;
assign  c[639:632]=8'h92;
assign  c[647:640]=8'h6c;
assign  c[655:648]=8'h70;
assign  c[663:656]=8'h48;
assign  c[671:664]=8'h50;
assign  c[679:672]=8'hfd;
assign  c[687:680]=8'hed;
assign  c[695:688]=8'hb9;
assign  c[703:696]=8'hda;
assign  c[711:704]=8'h5e;
assign  c[719:712]=8'h15;
assign  c[727:720]=8'h46;
assign  c[735:728]=8'h57;
assign  c[743:736]=8'ha7;
assign  c[751:744]=8'h8d;
assign  c[759:752]=8'h9d;
assign  c[767:760]=8'h84;
assign  c[775:768]=8'h90;
assign  c[783:776]=8'hd8;
assign  c[791:784]=8'hab;
assign  c[799:792]=8'h00;
assign  c[807:800]=8'h8c;
assign  c[815:808]=8'hbc;
assign  c[823:816]=8'hd3;
assign  c[831:824]=8'h0a;
assign  c[839:832]=8'hf7;
assign  c[847:840]=8'he4;
assign  c[855:848]=8'h58;
assign  c[863:856]=8'h05;
assign  c[871:864]=8'hb8;
assign  c[879:872]=8'hb3;
assign  c[887:880]=8'h45;
assign  c[895:888]=8'h06;
assign  c[903:896]=8'hd0;
assign  c[911:904]=8'h2c;
assign  c[919:912]=8'h1e;
assign  c[927:920]=8'h8f;
assign  c[935:928]=8'hca;
assign  c[943:936]=8'h3f;
assign  c[951:944]=8'h0f;
assign  c[959:952]=8'h02;
assign  c[967:960]=8'hc1;
assign  c[975:968]=8'haf;
assign  c[983:976]=8'hbd;
assign  c[991:984]=8'h03;
assign  c[999:992]=8'h01;
assign  c[1007:1000]=8'h13;
assign  c[1015:1008]=8'h8a;
assign  c[1023:1016]=8'h6b;
assign  c[1031:1024]=8'h3a;
assign  c[1039:1032]=8'h91;
assign  c[1047:1040]=8'h11;
assign  c[1055:1048]=8'h41;
assign  c[1063:1056]=8'h4f;
assign  c[1071:1064]=8'h67;
assign  c[1079:1072]=8'hdc;
assign  c[1087:1080]=8'hea;
assign  c[1095:1088]=8'h97;
assign  c[1103:1096]=8'hf2;
assign  c[1111:1104]=8'hcf;
assign  c[1119:1112]=8'hce;
assign  c[1127:1120]=8'hf0;
assign  c[1135:1128]=8'hb4;
assign  c[1143:1136]=8'he6;
assign  c[1151:1144]=8'h73;
assign  c[1159:1152]=8'h96;
assign  c[1167:1160]=8'hac;
assign  c[1175:1168]=8'h74;
assign  c[1183:1176]=8'h22;
assign  c[1191:1184]=8'he7;
assign  c[1199:1192]=8'had;
assign  c[1207:1200]=8'h35;
assign  c[1215:1208]=8'h85;
assign  c[1223:1216]=8'he2;
assign  c[1231:1224]=8'hf9;
assign  c[1239:1232]=8'h37;
assign  c[1247:1240]=8'he8;
assign  c[1255:1248]=8'h1c;
assign  c[1263:1256]=8'h75;
assign  c[1271:1264]=8'hdf;
assign  c[1279:1272]=8'h6e;
assign  c[1287:1280]=8'h47;
assign  c[1295:1288]=8'hf1;
assign  c[1303:1296]=8'h1a;
assign  c[1311:1304]=8'h71;
assign  c[1319:1312]=8'h1d;
assign  c[1327:1320]=8'h29;
assign  c[1335:1328]=8'hc5;
assign  c[1343:1336]=8'h89;
assign  c[1351:1344]=8'h6f;
assign  c[1359:1352]=8'hb7;
assign  c[1367:1360]=8'h62;
assign  c[1375:1368]=8'h0e;
assign  c[1383:1376]=8'haa;
assign  c[1391:1384]=8'h18;
assign  c[1399:1392]=8'hbe;
assign  c[1407:1400]=8'h1b;
assign  c[1415:1408]=8'hfc;
assign  c[1423:1416]=8'h56;
assign  c[1431:1424]=8'h3e;
assign  c[1439:1432]=8'h4b;
assign  c[1447:1440]=8'hc6;
assign  c[1455:1448]=8'hd2;
assign  c[1463:1456]=8'h79;
assign  c[1471:1464]=8'h20;
assign  c[1479:1472]=8'h9a;
assign  c[1487:1480]=8'hdb;
assign  c[1495:1488]=8'hc0;
assign  c[1503:1496]=8'hfe;
assign  c[1511:1504]=8'h78;
assign  c[1519:1512]=8'hcd;
assign  c[1527:1520]=8'h5a;
assign  c[1535:1528]=8'hf4;
assign  c[1543:1536]=8'h1f;
assign  c[1551:1544]=8'hdd;
assign  c[1559:1552]=8'ha8;
assign  c[1567:1560]=8'h33;
assign  c[1575:1568]=8'h88;
assign  c[1583:1576]=8'h07;
assign  c[1591:1584]=8'hc7;
assign  c[1599:1592]=8'h31;
assign  c[1607:1600]=8'hb1;
assign  c[1615:1608]=8'h12;
assign  c[1623:1616]=8'h10;
assign  c[1631:1624]=8'h59;
assign  c[1639:1632]=8'h27;
assign  c[1647:1640]=8'h80;
assign  c[1655:1648]=8'hec;
assign  c[1663:1656]=8'h5f;
assign  c[1671:1664]=8'h60;
assign  c[1679:1672]=8'h51;
assign  c[1687:1680]=8'h7f;
assign  c[1695:1688]=8'ha9;
assign  c[1703:1696]=8'h19;
assign  c[1711:1704]=8'hb5;
assign  c[1719:1712]=8'h4a;
assign  c[1727:1720]=8'h0d;
assign  c[1735:1728]=8'h2d;
assign  c[1743:1736]=8'he5;
assign  c[1751:1744]=8'h7a;
assign  c[1759:1752]=8'h9f;
assign  c[1767:1760]=8'h93;
assign  c[1775:1768]=8'hc9;
assign  c[1783:1776]=8'h9c;
assign  c[1791:1784]=8'hef;
assign  c[1799:1792]=8'ha0;
assign  c[1807:1800]=8'he0;
assign  c[1815:1808]=8'h3b;
assign  c[1823:1816]=8'h4d;
assign  c[1831:1824]=8'hae;
assign  c[1839:1832]=8'h2a;
assign  c[1847:1840]=8'hf5;
assign  c[1855:1848]=8'hb0;
assign  c[1863:1856]=8'hc8;
assign  c[1871:1864]=8'heb;
assign  c[1879:1872]=8'hbb;
assign  c[1887:1880]=8'h3c;
assign  c[1895:1888]=8'h83;
assign  c[1903:1896]=8'h53;
assign  c[1911:1904]=8'h99;
assign  c[1919:1912]=8'h61;
assign  c[1927:1920]=8'h17;
assign  c[1935:1928]=8'h2b;
assign  c[1943:1936]=8'h04;
assign  c[1951:1944]=8'h7e;
assign  c[1959:1952]=8'hba;
assign  c[1967:1960]=8'h77;
assign  c[1975:1968]=8'hd6;
assign  c[1983:1976]=8'h26;
assign  c[1991:1984]=8'he1;
assign  c[1999:1992]=8'h69;
assign  c[2007:2000]=8'h14;
assign  c[2015:2008]=8'h63;
assign  c[2023:2016]=8'h55;
assign  c[2031:2024]=8'h21;
assign  c[2039:2032]=8'h0c;
assign  c[2047:2040]=8'h7d;




wire[10:0] i0;
wire[10:0] i1;
wire[10:0] i2;
wire[10:0] i3;
wire[10:0] i4;
wire[10:0] i5;
wire[10:0] i6;
wire[10:0] i7;
wire[10:0] i8;
wire[10:0] i9;
wire[10:0] i10;
wire[10:0] i11;
wire[10:0] i12;
wire[10:0] i13;
wire[10:0] i14;
wire[10:0] i15;

assign i0 = 'd128* stateIn[7:4] + 'd8*stateIn[3:0];
assign stateOut[7:0] = c[ i0 +: 8];

assign i1 = 'd128* stateIn[15:12] + 'd8*stateIn[11:8];
assign stateOut[15:8] = c[ i1 +: 8];

assign i2 = 'd128* stateIn[23:20] + 'd8*stateIn[19:16];
assign stateOut[23:16] = c[ i2 +: 8];

assign i3 = 'd128* stateIn[31:28] + 'd8*stateIn[27:24];
assign stateOut[31:24] = c[ i3 +: 8];

assign i4 = 'd128* stateIn[39:36] + 'd8*stateIn[35:32];
assign stateOut[39:32] = c[ i4 +: 8];

assign i5 = 'd128* stateIn[47:44] + 'd8*stateIn[43:40];
assign stateOut[47:40] = c[ i5 +: 8];

assign i6 = 'd128* stateIn[55:52] + 'd8*stateIn[51:48] ;
assign stateOut[55:48] = c[ i6 +: 8 ];

assign i7 = 'd128* stateIn[63:60] + 'd8*stateIn[59:56];
assign stateOut[63:56] = c[ i7 +: 8];

assign i8 = 'd128* stateIn[71:68] + 'd8*stateIn[67:64];
assign stateOut[71:64] = c[ i8 +: 8];

assign i9 = 'd128* stateIn[79:76] + 'd8*stateIn[75:72];
assign stateOut[79:72] = c[ i9 +: 8];

assign i10 = 'd128* stateIn[87:84] + 'd8*stateIn[83:80];
assign stateOut[87:80] = c[ i10 +: 8];

assign i11 = 'd128* stateIn[95:92] + 'd8*stateIn[91:88];
assign stateOut[95:88] = c[ i11 +: 8];

assign i12 = 'd128* stateIn[103:100] + 'd8*stateIn[99:96];
assign stateOut[103:96] = c[ i12 +: 8];

assign i13 = 'd128* stateIn[111:108] + 'd8*stateIn[107:104];
assign stateOut[111:104] = c[ i13 +: 8];

assign i14 = 'd128* stateIn[119:116] + 'd8*stateIn[115:112];
assign stateOut[119:112] = c[ i14 +: 8];

assign i15 = 'd128* stateIn[127:124] + 'd8*stateIn[123:120];
assign stateOut[127:120] = c[ i15 +: 8];

endmodule
 
